`ifndef INSTRUCTIONS_H
`define INSTRUCTIONS_H

`include "instructions/ora.svh"

`endif