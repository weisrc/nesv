`ifndef MATRIX_H
`define MATRIX_H

`include "matrix/0.sv"
`include "matrix/4.sv"
`include "matrix/8.sv"
`include "matrix/A.sv"
`include "matrix/C.sv"
`include "matrix/1259D.sv"
`include "matrix/6E.sv"

`endif
