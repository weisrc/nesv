`include "../common.sv"
`include "../actions.sv"

function void column_6(inout state_t state);
  case (state.op[7:4])

    'h0: begin
    end
    'h1: begin
    end
    'h2: begin
    end
    'h3: begin
    end
    'h4: begin
    end
    'h5: begin
    end
    'h6: begin
    end
    'h7: begin
    end
    'h8: begin
    end
    'h9: begin
    end
    'hA: begin
    end
    'hB: begin
    end
    'hC: begin
    end
    'hD: begin
    end
    'hE: begin
    end
    'hF: begin
    end

  endcase
endfunction
