`ifndef MATRIX_H
`define MATRIX_H

`include "matrix/0.sv"
`include "matrix/1.sv"
`include "matrix/2.sv"
`include "matrix/3.sv"
`include "matrix/4.sv"
`include "matrix/5.sv"
`include "matrix/6.sv"
`include "matrix/7.sv"
`include "matrix/8.sv"
`include "matrix/9.sv"
`include "matrix/A.sv"
`include "matrix/B.sv"
`include "matrix/C.sv"
`include "matrix/D.sv"
`include "matrix/E.sv"
`include "matrix/F.sv"

`endif
