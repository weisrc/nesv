`include "../common.sv"

`ifndef BRANCHING_H
`define BRANCHING_H

`endif