`ifndef COLUMNS_H
`define COLUMNS_H

`include "columns/0.svh"
`include "columns/1.svh"
`include "columns/2.svh"
`include "columns/3.svh"
`include "columns/4.svh"
`include "columns/5.svh"
`include "columns/6.svh"
`include "columns/7.svh"
`include "columns/8.svh"
`include "columns/9.svh"
`include "columns/A.svh"
`include "columns/B.svh"
`include "columns/C.svh"
`include "columns/D.svh"
`include "columns/E.svh"
`include "columns/F.svh"

`endif