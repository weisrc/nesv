`ifndef ACTIONS_H
`define ACTIONS_H

`include "actions/bitwise.sv"
`include "actions/modes.sv"
`include "actions/memory.sv"

`endif