`include "../common.sv"
`include "../actions.sv"

function void column_A(inout state_t state); case (state.op[7:4])

4'h0: begin end
4'h1: begin end
4'h2: begin end
4'h3: begin end
4'h4: begin end
4'h5: begin end
4'h6: begin end
4'h7: begin end
4'h8: begin end
4'h9: begin end
4'hA: begin end
4'hB: begin end
4'hC: begin end
4'hD: begin end
4'hE: begin end
4'hF: begin end

endcase endfunction