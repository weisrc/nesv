`ifndef COLUMNS_H
`define COLUMNS_H

`include "columns/0.sv"
`include "columns/1.sv"
`include "columns/2.sv"
`include "columns/3.sv"
`include "columns/4.sv"
`include "columns/5.sv"
`include "columns/6.sv"
`include "columns/7.sv"
`include "columns/8.sv"
`include "columns/9.sv"
`include "columns/A.sv"
`include "columns/B.sv"
`include "columns/C.sv"
`include "columns/D.sv"
`include "columns/E.sv"
`include "columns/F.sv"

`endif
