`ifndef ACTIONS_H
`define ACTIONS_H

`include "actions/bitwise.sv"
`include "actions/addressing.sv"
`include "actions/memory.sv"
`include "actions/status.sv"
`include "actions/arithmetic.sv"

`endif