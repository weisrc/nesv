`ifndef MODES_H
`define MODES_H

`include "modes/read_ind_x.svh"

`endif