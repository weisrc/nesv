`ifndef ACTIONS_H
`define ACTIONS_H

`include "actions/bitwise.sv"
`include "actions/branching.sv"
`include "actions/addressing.sv"
`include "actions/memory.sv"
`include "actions/status.sv"
`include "actions/arithmetic.sv"
`include "actions/shifting.sv"
`include "actions/stack.sv"
`include "actions/compare.sv"
`include "actions/transfer.sv"

`endif
